package router_test_pkg;

        import uvm_pkg::*;

        `include "uvm_macros.svh"

        `include "src_config.sv"
        `include "dst_config.sv"
        `include "env_config.sv"

        `include "src_xtn.sv"
        `include "src_seq.sv"
        `include "src_seqr.sv"
        `include "src_mon.sv"
        `include "src_drv.sv"
        `include "src_agt.sv"
        `include "src_agt_top.sv"

        `include "dst_xtn.sv"
        `include "dst_sequence.sv"
        `include "dst_sequencer.sv"
        `include "dst_monitor.sv"
        `include "dst_driver.sv"
        `include "dst_agt.sv"
        `include "dst_agt_top.sv"

        `include "router_virtual_sequencer.sv"
        `include "router_virtual_sequence.sv"
        `include "scoreboard.sv"
        `include "router_env.sv"
        `include "router_test.sv"

endpackage
